0010001000000011011001011010010000000000000000001100000000000000000000000000011000000000000000000000000000000000010011
0010001000000011011011010010010000000000000000000001000000000000000000000000000010000000000000000000000000000000110001
0110001000000011101110110100010000000000000000011111100000000000000000000000111111000000000000000000000000000000000000
0110001000000101101001110111010000000000000000000001000000000000000000000000000010000000000000000000000000000000000000
