000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100
000010001000000011011000111110010000000000000000000000000000001111110000000000000000000000000000000100000000000000000000000000011100000000000000000000000000000111001000100000000000000000000000000000000000000000000000000000010100000000000000000000000000000000010000000000000000000000000000010100000000000000000000000000000101
000010001000000011011001011010010000000000000000000000000000001111110000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000011001000100000000000000001010000000000000000000000000000000000110010000000000000000000000000000101000000000000000000000000000000010100000000000000000000000000000101
000110001000000011011011010010010000000000000000000000000000001111110000000000000000000000000011001000000000000000000000000000000100000000000000000000000000000001001000100000000000111111110000000000000000000000000000000111110100000000000000000000000000000000010000000000000000000000110010000000000000000000000000000000000001
000110001000000011101110110100010000000000000000000000000000001111110000000000000000000000011111010000000000000000000000000000000001000000000000000000000000000000011000100000001101010100001111000000000000000000000000000000001010000000000000000000000000000000010000000000000000000000011111010000000000000000000000000000000001
