000000000000000111000010001000000011011000111110010000000000000000111000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000
000000000000000001100010001000000011011001011010010000000000000000001100000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000000000000000000000000110001000000000000000000000000000000000000000000000000100010001000000000000000010100000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000
010000110001010001111110001000000000001111111100000000000110001010001111100000000000001100010100011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010001000000011011011010010010000000000000000110010000000000000000000000001100100000000000000000000000000000000000000
010000000000111110101010001000000011010101000011110000000000000111110101000000000000000000001111101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111010001000000011101110110100010000000000000000011111100000000000000000000000111111000000000000000000000000000000000000
